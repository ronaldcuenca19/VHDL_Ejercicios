----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    11:38:14 05/23/2022 
-- Design Name: 
-- Module Name:    ejercicio2_Suma - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity ejercicio2_Suma is
Port ( 
           A : in bit_vector (0 to 1);
			  B : in bit_vector (0 to 1);
			  suma : out bit_vector (0 to 1));
end ejercicio2_Suma;

architecture Behavioral of ejercicio2_Suma is

begin


end Behavioral;

